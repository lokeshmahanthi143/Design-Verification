module ;
endmodule 

