module;
endmodule 
